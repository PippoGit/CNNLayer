library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.cnn_types.all;

entity CNNFilterRom is
  port (
    filter_3x3 : out cnn_matrix_t(0 to 2, 0 to 2);
    filter_4x4 : out cnn_matrix_t(0 to 3, 0 to 3);
    filter_6x6 : out cnn_matrix_t(0 to 5, 0 to 5)
  );
end CNNFilterRom;

architecture CNNFilterRom_Arch of CNNFilterRom is
begin
  filter_3x3 <= (
     ("00000001", "00000000", "00000001"),
     ("00000000", "00000001", "00000000"),
     ("00000001", "00000000", "00000001") 
  );

  filter_4x4 <= (
     ("00000000", "00000000", "00000000", "00000000"),
     ("00000000", "00000000", "00000000", "00000000"),
     ("00000000", "00000000", "00000000", "00000000"),
     ("00000000", "00000000", "00000000", "00000000")  
  );

  filter_6x6 <= (
    ("00000000", "00000000", "00000000", "00000000", "00000000", "00000000"),
    ("00000000", "00000000", "00000000", "00000000", "00000000", "00000000"),
    ("00000000", "00000000", "00000000", "00000000", "00000000", "00000000"),
    ("00000000", "00000000", "00000000", "00000000", "00000000", "00000000"),
    ("00000000", "00000000", "00000000", "00000000", "00000000", "00000000"),
    ("00000000", "00000000", "00000000", "00000000", "00000000", "00000000")
  );
end CNNFilterRom_Arch;
